sebastien lauret    fqd1235             26 parc de la berengere                           saint cloud         france                      �       p�@{       sebastien lauret    fqd1235             26 parc de la berengere                           saint cloud         france                      �       p�@{       