seb       lau       123D                26 parc de la berengere                           saint cloud         frnace                      �       p�@       